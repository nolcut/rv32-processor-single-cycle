module beaver32rv (input wire clk;);
    
endmodule